`timescale 20ns/20ns
module gDMA ();
    
endmodule